package com.disb;

import javax.persistence.*;
import java.io.Serializable;
import java.util.Objects;

/*
@Entity
@Table(name = "ahli")
@Cache(usage = CacheConcurrencyStrategy.NONSTRICT_READ_WRITE)
public class Ahli implements Serializable {

	@Id
    @GeneratedValue(strategy = GenerationType.AUTO)
    private Long id;

    @Column(name = "kp")
    private String kp;
    
    @Column(name = "nama")
    private String nama;
    
    @Column(name = "tel")
    private String tel;
    
    @Column(name = "emel")
    private String emel;

    @Column(name = "alamat")
    private String alamat;

    public Long getId() {
        return id;
    }

    public void setId(Long id) {
        this.id = id;
    }

    public String getKp() {
        return kp;
    }
    
    public void setKp(String kp) {
        this.kp = kp;
    }

    public String getNama() {
        return nama;
    }
    
    public void setNama(String nama) {
        this.nama = nama;
    }

    public String getTel() {
        return tel;
    }
    
    public void setTel(String tel) {
        this.tel = tel;
    }

    public String getEmel() {
        return emel;
    }
    
    public void setEmel(String emel) {
        this.emel = emel;
    }

    public String getAlamat() {
        return alamat;
    }
    
    public void setAlamat(String alamat) {
        this.alamat = alamat;
    }

    @Override
    public String toString() {
        return "Ahli{" +
            "id=" + id +
            ", kp='" + kp + "'" +
            ", nama='" + nama + "'" +
            ", tel='" + tel + "'" +
            ", emel='" + emel + "'" +
            ", alamat='" + alamat + "'" +
            '}';
    }

}
*/

